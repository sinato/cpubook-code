module and_mod(
    input x,
    input y,
    output z
);
    assign z = x & y;
endmodule